    //
	// USER LOGIC
    //

    import hash_table::*;
    import linked_list::*;
    
    dlm_1t2n1c8p inst_user_logic_dlm (

        .axi_ctrl_awvalid(axi_ctrl_user.awvalid),
        .axi_ctrl_awready(axi_ctrl_user.awready),
        .axi_ctrl_awaddr(axi_ctrl_user.awaddr),
        .axi_ctrl_awprot(),
        .axi_ctrl_wvalid(axi_ctrl_user.wvalid),
        .axi_ctrl_wready(axi_ctrl_user.wready),
        .axi_ctrl_wdata(axi_ctrl_user.wdata),
        .axi_ctrl_wstrb(axi_ctrl_user.wstrb),
        .axi_ctrl_arvalid(axi_ctrl_user.arvalid),
        .axi_ctrl_arready(axi_ctrl_user.arready),
        .axi_ctrl_araddr(axi_ctrl_user.araddr),
        .axi_ctrl_arprot(),
        .axi_ctrl_rvalid(axi_ctrl_user.rvalid),
        .axi_ctrl_rready(axi_ctrl_user.rready),
        .axi_ctrl_rdata(axi_ctrl_user.rdata),
        .axi_ctrl_rresp(axi_ctrl_user.rresp),
        .axi_ctrl_bvalid(axi_ctrl_user.bvalid),
        .axi_ctrl_bready(axi_ctrl_user.bready),
        .axi_ctrl_bresp(axi_ctrl_user.bresp),

        .hostd_bpss_rd_req_data(bpss_rd_req.data),
        .hostd_bpss_rd_req_valid(bpss_rd_req.valid),
        .hostd_bpss_rd_req_ready(bpss_rd_req.ready),
        .hostd_bpss_wr_req_data(bpss_wr_req.data),
        .hostd_bpss_wr_req_valid(bpss_wr_req.valid),
        .hostd_bpss_wr_req_ready(bpss_wr_req.ready),
        .hostd_bpss_rd_done_data(bpss_rd_done.data),
        .hostd_bpss_rd_done_valid(bpss_rd_done.valid),
        .hostd_bpss_rd_done_ready(),
        .hostd_bpss_wr_done_data(bpss_wr_done.data),
        .hostd_bpss_wr_done_valid(bpss_wr_done.valid),
        .hostd_bpss_wr_done_ready(),

        .hostd_axis_host_sink_tdata(axis_host_sink_mux[0].tdata),
        .hostd_axis_host_sink_tkeep(axis_host_sink_mux[0].tkeep),
        .hostd_axis_host_sink_tdest(axis_host_sink_mux[0].tid),
        .hostd_axis_host_sink_tlast(axis_host_sink_mux[0].tlast),
        .hostd_axis_host_sink_tvalid(axis_host_sink_mux[0].tvalid),
        .hostd_axis_host_sink_tready(axis_host_sink_mux[0].tready),
        .hostd_axis_host_src_tdata(axis_host_src_mux[0].tdata),
        .hostd_axis_host_src_tkeep(axis_host_src_mux[0].tkeep),
        .hostd_axis_host_src_tdest(axis_host_src_mux[0].tid),
        .hostd_axis_host_src_tlast(axis_host_src_mux[0].tlast),
        .hostd_axis_host_src_tvalid(axis_host_src_mux[0].tvalid),
        .hostd_axis_host_src_tready(axis_host_src_mux[0].tready),

            .axi_mem_0_awvalid(axi_mem_0_awvalid),
            .axi_mem_0_awready(axi_mem_0_awready),
            .axi_mem_0_awaddr(axi_mem_0_awaddr),
            .axi_mem_0_awid(axi_mem_0_awid),
            .axi_mem_0_awlen(axi_mem_0_awlen),
            .axi_mem_0_awsize(axi_mem_0_awsize),
            .axi_mem_0_awburst(axi_mem_0_awburst),

            .axi_mem_0_wvalid(axi_mem_0_wvalid),
            .axi_mem_0_wready(axi_mem_0_wready),
            .axi_mem_0_wdata(axi_mem_0_wdata),
            .axi_mem_0_wstrb(axi_mem_0_wstrb),
            .axi_mem_0_wlast(axi_mem_0_wlast),
            .axi_mem_0_bvalid(axi_mem_0_bvalid),
            .axi_mem_0_bready(axi_mem_0_bready),
            .axi_mem_0_bid(axi_mem_0_bid),
            .axi_mem_0_bresp(axi_mem_0_bresp),

            .axi_mem_0_arvalid(axi_mem_0_arvalid),
            .axi_mem_0_arready(axi_mem_0_arready),
            .axi_mem_0_araddr(axi_mem_0_araddr),
            .axi_mem_0_arid(axi_mem_0_arid),
            .axi_mem_0_arlen(axi_mem_0_arlen),
            .axi_mem_0_arsize(axi_mem_0_arsize),
            .axi_mem_0_arburst(axi_mem_0_arburst),

            .axi_mem_0_rvalid(axi_mem_0_rvalid),
            .axi_mem_0_rready(axi_mem_0_rready),
            .axi_mem_0_rdata(axi_mem_0_rdata),
            .axi_mem_0_rid(axi_mem_0_rid),
            .axi_mem_0_rresp(axi_mem_0_rresp),
            .axi_mem_0_rlast(axi_mem_0_rlast),

            .axi_mem_1_awvalid(axi_mem_1_awvalid),
            .axi_mem_1_awready(axi_mem_1_awready),
            .axi_mem_1_awaddr(axi_mem_1_awaddr),
            .axi_mem_1_awid(axi_mem_1_awid),
            .axi_mem_1_awlen(axi_mem_1_awlen),
            .axi_mem_1_awsize(axi_mem_1_awsize),
            .axi_mem_1_awburst(axi_mem_1_awburst),

            .axi_mem_1_wvalid(axi_mem_1_wvalid),
            .axi_mem_1_wready(axi_mem_1_wready),
            .axi_mem_1_wdata(axi_mem_1_wdata),
            .axi_mem_1_wstrb(axi_mem_1_wstrb),
            .axi_mem_1_wlast(axi_mem_1_wlast),
            .axi_mem_1_bvalid(axi_mem_1_bvalid),
            .axi_mem_1_bready(axi_mem_1_bready),
            .axi_mem_1_bid(axi_mem_1_bid),
            .axi_mem_1_bresp(axi_mem_1_bresp),

            .axi_mem_1_arvalid(axi_mem_1_arvalid),
            .axi_mem_1_arready(axi_mem_1_arready),
            .axi_mem_1_araddr(axi_mem_1_araddr),
            .axi_mem_1_arid(axi_mem_1_arid),
            .axi_mem_1_arlen(axi_mem_1_arlen),
            .axi_mem_1_arsize(axi_mem_1_arsize),
            .axi_mem_1_arburst(axi_mem_1_arburst),

            .axi_mem_1_rvalid(axi_mem_1_rvalid),
            .axi_mem_1_rready(axi_mem_1_rready),
            .axi_mem_1_rdata(axi_mem_1_rdata),
            .axi_mem_1_rid(axi_mem_1_rid),
            .axi_mem_1_rresp(axi_mem_1_rresp),
            .axi_mem_1_rlast(axi_mem_1_rlast),

            .axi_mem_2_awvalid(axi_mem_2_awvalid),
            .axi_mem_2_awready(axi_mem_2_awready),
            .axi_mem_2_awaddr(axi_mem_2_awaddr),
            .axi_mem_2_awid(axi_mem_2_awid),
            .axi_mem_2_awlen(axi_mem_2_awlen),
            .axi_mem_2_awsize(axi_mem_2_awsize),
            .axi_mem_2_awburst(axi_mem_2_awburst),

            .axi_mem_2_wvalid(axi_mem_2_wvalid),
            .axi_mem_2_wready(axi_mem_2_wready),
            .axi_mem_2_wdata(axi_mem_2_wdata),
            .axi_mem_2_wstrb(axi_mem_2_wstrb),
            .axi_mem_2_wlast(axi_mem_2_wlast),
            .axi_mem_2_bvalid(axi_mem_2_bvalid),
            .axi_mem_2_bready(axi_mem_2_bready),
            .axi_mem_2_bid(axi_mem_2_bid),
            .axi_mem_2_bresp(axi_mem_2_bresp),

            .axi_mem_2_arvalid(axi_mem_2_arvalid),
            .axi_mem_2_arready(axi_mem_2_arready),
            .axi_mem_2_araddr(axi_mem_2_araddr),
            .axi_mem_2_arid(axi_mem_2_arid),
            .axi_mem_2_arlen(axi_mem_2_arlen),
            .axi_mem_2_arsize(axi_mem_2_arsize),
            .axi_mem_2_arburst(axi_mem_2_arburst),

            .axi_mem_2_rvalid(axi_mem_2_rvalid),
            .axi_mem_2_rready(axi_mem_2_rready),
            .axi_mem_2_rdata(axi_mem_2_rdata),
            .axi_mem_2_rid(axi_mem_2_rid),
            .axi_mem_2_rresp(axi_mem_2_rresp),
            .axi_mem_2_rlast(axi_mem_2_rlast),

            .axi_mem_3_awvalid(axi_mem_3_awvalid),
            .axi_mem_3_awready(axi_mem_3_awready),
            .axi_mem_3_awaddr(axi_mem_3_awaddr),
            .axi_mem_3_awid(axi_mem_3_awid),
            .axi_mem_3_awlen(axi_mem_3_awlen),
            .axi_mem_3_awsize(axi_mem_3_awsize),
            .axi_mem_3_awburst(axi_mem_3_awburst),

            .axi_mem_3_wvalid(axi_mem_3_wvalid),
            .axi_mem_3_wready(axi_mem_3_wready),
            .axi_mem_3_wdata(axi_mem_3_wdata),
            .axi_mem_3_wstrb(axi_mem_3_wstrb),
            .axi_mem_3_wlast(axi_mem_3_wlast),
            .axi_mem_3_bvalid(axi_mem_3_bvalid),
            .axi_mem_3_bready(axi_mem_3_bready),
            .axi_mem_3_bid(axi_mem_3_bid),
            .axi_mem_3_bresp(axi_mem_3_bresp),

            .axi_mem_3_arvalid(axi_mem_3_arvalid),
            .axi_mem_3_arready(axi_mem_3_arready),
            .axi_mem_3_araddr(axi_mem_3_araddr),
            .axi_mem_3_arid(axi_mem_3_arid),
            .axi_mem_3_arlen(axi_mem_3_arlen),
            .axi_mem_3_arsize(axi_mem_3_arsize),
            .axi_mem_3_arburst(axi_mem_3_arburst),

            .axi_mem_3_rvalid(axi_mem_3_rvalid),
            .axi_mem_3_rready(axi_mem_3_rready),
            .axi_mem_3_rdata(axi_mem_3_rdata),
            .axi_mem_3_rid(axi_mem_3_rid),
            .axi_mem_3_rresp(axi_mem_3_rresp),
            .axi_mem_3_rlast(axi_mem_3_rlast),
            
        .rdma_0_rd_req_data(rdma_0_rd_req.data),
        .rdma_0_rd_req_valid(rdma_0_rd_req.valid),
        .rdma_0_rd_req_ready(rdma_0_rd_req.ready),
        .rdma_0_wr_req_data(rdma_0_wr_req_mux.data),
        .rdma_0_wr_req_valid(rdma_0_wr_req_mux.valid),
        .rdma_0_wr_req_ready(rdma_0_wr_req_mux.ready),
        .rdma_0_sq_data(rdma_0_sq.data),
        .rdma_0_sq_valid(rdma_0_sq.valid),
        .rdma_0_sq_ready(rdma_0_sq.ready),
        .rdma_0_ack_data(rdma_0_ack.data),
        .rdma_0_ack_valid(rdma_0_ack.valid),
        .rdma_0_ack_ready(rdma_0_ack.ready),
        .rdma_0_axis_sink_tdata(axis_rdma_0_sink_mux.tdata),
        .rdma_0_axis_sink_tkeep(axis_rdma_0_sink_mux.tkeep),
        // .rdma_0_axis_sink_tid(axis_rdma_0_sink_mux.tid),
        .rdma_0_axis_sink_tlast(axis_rdma_0_sink_mux.tlast),
        .rdma_0_axis_sink_tvalid(axis_rdma_0_sink_mux.tvalid),
        .rdma_0_axis_sink_tready(axis_rdma_0_sink_mux.tready),
        .rdma_0_axis_src_tdata(axis_rdma_0_src.tdata),
        .rdma_0_axis_src_tkeep(axis_rdma_0_src.tkeep),
        // .rdma_0_axis_src_tid(axis_rdma_0_src.tid),
        .rdma_0_axis_src_tlast(axis_rdma_0_src.tlast),
        .rdma_0_axis_src_tvalid(axis_rdma_0_src.tvalid),
        .rdma_0_axis_src_tready(axis_rdma_0_src.tready),

        .resetn(aresetn),
        .clk(aclk)
	);